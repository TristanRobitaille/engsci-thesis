`ifndef _cim_svh_
`define _cim_svh_

/*----- ENUM -----*/
    typedef enum logic [2:0] {
        CIM_IDLE,
        CIM_RESET,
        CIM_PATCH_LOAD,
        CIM_INFERENCE_RUNNING,
        CIM_INVALID,
        CIM_NUM_STATES
    } CIM_STATE_T;

    typedef enum logic [5:0] {
        CLASS_TOKEN_CONCAT_STEP,
        POS_EMB_STEP,
        ENC_LAYERNORM_1_1ST_HALF_STEP,
        ENC_LAYERNORM_1_2ND_HALF_STEP,
        ENC_LAYERNORM_2_1ST_HALF_STEP,
        ENC_LAYERNORM_2_2ND_HALF_STEP,
        ENC_LAYERNORM_3_1ST_HALF_STEP,
        ENC_LAYERNORM_3_2ND_HALF_STEP,
        POST_LAYERNORM_TRANSPOSE_STEP,
        ENC_MHSA_DENSE_STEP,
        ENC_MHSA_Q_TRANSPOSE_STEP,
        ENC_MHSA_K_TRANSPOSE_STEP,
        ENC_MHSA_QK_T_STEP,
        ENC_MHSA_PRE_SOFTMAX_TRANSPOSE_STEP,
        ENC_MHSA_SOFTMAX_STEP,
        ENC_MHSA_MULT_V_STEP,
        ENC_POST_MHSA_TRANSPOSE_STEP,
        ENC_POST_MHSA_DENSE_AND_INPUT_SUM_STEP,
        ENC_PRE_MLP_TRANSPOSE_STEP,
        MLP_DENSE_1_STEP,
        ENC_POST_DENSE_1_TRANSPOSE_STEP,
        MLP_DENSE_2_AND_SUM_STEP,
        MLP_HEAD_PRE_DENSE_1_TRANSPOSE_STEP,
        MLP_HEAD_DENSE_1_STEP,
        MLP_HEAD_PRE_DENSE_2_TRANSPOSE_STEP,
        MLP_HEAD_DENSE_2_STEP,
        MLP_HEAD_PRE_SOFTMAX_TRANSPOSE_STEP,
        MLP_HEAD_SOFTMAX_STEP,
        POST_SOFTMAX_DIVIDE_STEP,
        POST_SOFTMAX_AVERAGING_STEP,
        RETIRE_SOFTMAX_STEP,
        INFERENCE_COMPLETE,
        INVALID_INF_STEP
    } INFERENCE_STEP_T;

`endif
