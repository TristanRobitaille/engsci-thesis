`ifndef _master_init_sv_
`define _master_init_sv_

`include "master.svh"

const BroadcastOpInfo_t broadcast_ops[25] = '{ 
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+3*(NUM_PATCHES+1)),  /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+3*(NUM_PATCHES+1)),  /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+NUM_PATCHES+1),      /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*(EMB_DEPTH+NUM_PATCHES+1)),    /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+NUM_PATCHES+1),      /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*len*/ $clog2(NUM_CIMS+1)'(NUM_HEADS),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(3*EMB_DEPTH+NUM_PATCHES+1),      /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(3*EMB_DEPTH+2*(NUM_PATCHES+1)),  /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*(EMB_DEPTH+NUM_PATCHES+1)),    /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ NOP,                        /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*len*/ $clog2(NUM_CIMS+1)'(0),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*num_cim*/ $clog2(NUM_CIMS+1)'(0)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*(EMB_DEPTH+NUM_PATCHES+1)),    /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+NUM_PATCHES+1),      /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH+NUM_PATCHES+1),      /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*len*/ $clog2(NUM_CIMS+1)'(NUM_PATCHES+1), /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(4*EMB_DEPTH+NUM_PATCHES+1),      /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(4*EMB_DEPTH+NUM_PATCHES+1),      /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1+EMB_DEPTH),        /*len*/ $clog2(NUM_CIMS+1)'(1),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(MLP_DIM)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*len*/ $clog2(NUM_CIMS+1)'(MLP_DIM),       /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(NUM_PATCHES+1),                  /*num_cim*/ $clog2(NUM_CIMS+1)'(1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(3*EMB_DEPTH+NUM_PATCHES+2),      /*len*/ $clog2(NUM_CIMS+1)'(1),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_CIMS)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(EMB_DEPTH),                      /*num_cim*/ $clog2(NUM_CIMS+1)'(1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(EMB_DEPTH),                      /*len*/ $clog2(NUM_CIMS+1)'(1),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*num_cim*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*len*/ $clog2(NUM_CIMS+1)'(EMB_DEPTH),     /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(EMB_DEPTH),                      /*num_cim*/ $clog2(NUM_CIMS+1)'(1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH),                    /*len*/ $clog2(NUM_CIMS+1)'(1),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(0),                              /*num_cim*/ $clog2(NUM_CIMS+1)'(MLP_DIM)},
    {/*op*/ DENSE_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(MLP_DIM),                        /*len*/ $clog2(NUM_CIMS+1)'(MLP_DIM),       /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(EMB_DEPTH),                      /*num_cim*/ $clog2(NUM_CIMS+1)'(1)},
    {/*op*/ TRANS_BROADCAST_START_OP,   /*tx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(2*EMB_DEPTH),                    /*len*/ $clog2(NUM_CIMS+1)'(1),             /*rx_addr*/ $clog2(TEMP_RES_STORAGE_SIZE_CIM)'(MLP_DIM),                        /*num_cim*/ $clog2(NUM_CIMS+1)'(NUM_SLEEP_STAGES)}
};

`endif
