`ifndef _cim_centralized_vh_
`define _cim_centralized_vh_

import Defines::*;

module cim_centralized #()(
    input wire clk,
    SoCInterface soc_ctrl_i,

    // ----- Memory ---- //
    output MemoryInterface.input_write  param_write_tb_i,
    output MemoryInterface.input_write int_res_write_tb_i
);
    // ----- INSTANTIATION ----- //
    // Counters
    CounterInterface #(.WIDTH(4)) cnt_4b_i ();
    CounterInterface #(.WIDTH(7)) cnt_7b_i ();
    CounterInterface #(.WIDTH(9)) cnt_9b_i ();
    counter #(.WIDTH(4), .MODE(LEVEL_TRIGGERED)) cnt_4b_u (.clk(clk), .sig(cnt_4b_i));
    counter #(.WIDTH(7), .MODE(LEVEL_TRIGGERED)) cnt_7b_u (.clk(clk), .sig(cnt_7b_i));
    counter #(.WIDTH(9), .MODE(LEVEL_TRIGGERED)) cnt_9b_u (.clk(clk), .sig(cnt_9b_i));

    // Memory
    MemoryInterface #(CompFx_t, ParamAddr_t, FxFormatParams_t) param_write_i ();
    MemoryInterface #(CompFx_t, ParamAddr_t, FxFormatParams_t) param_read_i ();
    MemoryInterface #(CompFx_t, ParamAddr_t, FxFormatParams_t) param_read_mac_i ();
    MemoryInterface #(CompFx_t, ParamAddr_t, FxFormatParams_t) param_read_cim_i ();
    MemoryInterface #(CompFx_t, ParamAddr_t, FxFormatParams_t) param_read_ln_i ();

    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_read_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_write_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_read_cim_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_read_mac_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_read_ln_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_write_cim_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) int_res_write_ln_i ();

    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) mac_casts_i ();
    MemoryInterface #(CompFx_t, IntResAddr_t, FxFormatIntRes_t) ln_casts_i ();

    params_mem params_u   (.clk, .rst_n, .write(param_write_tb_i),.read(param_read_i)); // Only testbench writes to params
    int_res_mem int_res_u (.clk, .rst_n, .write(int_res_write_i), .read(int_res_read_i));

    // Compute
    ComputeIPInterface add_io();
    ComputeIPInterface add_io_cim();
    ComputeIPInterface add_io_exp();
    ComputeIPInterface add_io_mac();
    ComputeIPInterface add_io_ln();
    ComputeIPInterface mult_io();
    ComputeIPInterface mult_io_exp();
    ComputeIPInterface mult_io_mac();
    ComputeIPInterface mult_io_ln();
    ComputeIPInterface div_io();
    ComputeIPInterface div_io_mac();
    ComputeIPInterface div_io_ln();
    ComputeIPInterface exp_io();
    ComputeIPInterface exp_io_mac();
    ComputeIPInterface sqrt_io();
    ComputeIPInterface mac_io();
    ComputeIPInterface mac_io_extra();
    ComputeIPInterface ln_io();
    ComputeIPInterface ln_io_extra();

    adder add       (.clk, .rst_n, .io(add_io));
    multiplier mult (.clk, .rst_n, .io(mult_io));
    divider div     (.clk, .rst_n, .io(div_io));
    exp exp         (.clk, .rst_n, .io(exp_io), .adder_io(add_io_exp), .mult_io(mult_io_exp));
    sqrt sqrt       (.clk, .rst_n, .io(sqrt_io));
    mac mac         (.clk, .rst_n, .io(mac_io), .io_extra(mac_io_extra),
                     .casts(mac_casts_i), .param_read(param_read_mac_i), .int_res_read(int_res_read_mac_i),
                     .add_io(add_io_mac), .mult_io(mult_io_mac), .div_io(div_io_mac), .exp_io(exp_io_mac));
    layernorm layernorm (.clk, .rst_n, .io(ln_io), .io_extra(ln_io_extra), .add_io(add_io_ln), .mult_io(mult_io_ln), .div_io(div_io_ln), .sqrt_io,
                         .casts(ln_casts_i), .param_read(param_read_ln_i), .int_res_read(int_res_read_ln_i), .int_res_write(int_res_write_ln_i));

    // ----- GLOBAL SIGNALS ----- //
    logic rst_n;
    logic [1:0] delay_line_2b;
    State_t cim_state;
    InferenceStep_t current_inf_step;

    // ----- CONSTANTS -----//
    assign rst_n = soc_ctrl_i.rst_n;

    // ----- FSM ----- //
    always_ff @ (posedge clk) begin : main_fsm
        if (~rst_n) begin
            reset();
        end else begin
            unique case (cim_state)
                IDLE_CIM: begin
                    current_inf_step <= PATCH_PROJ_STEP;
                    if (soc_ctrl_i.start_eeg_load) cim_state <= EEG_LOAD;
                    if (soc_ctrl_i.new_sleep_epoch) cim_state <= INFERENCE_RUNNING;
                end
                EEG_LOAD: begin
                    if (soc_ctrl_i.new_sleep_epoch) cim_state <= INFERENCE_RUNNING;
                end
                INFERENCE_RUNNING: begin
                    if (current_inf_step == ENC_LAYERNORM_1_2ND_HALF_STEP) begin
                        cim_state <= IDLE_CIM;
                        soc_ctrl_i.inference_complete <= 1'b1;
                    end
                end
                INVALID_CIM: begin
                    cim_state <= IDLE_CIM;
                end
                default: begin
                    cim_state <= IDLE_CIM;
                end
            endcase
        end
    end

    always_ff @ (posedge clk) begin : inference_fsm
        set_default_values();
        if (cim_state == EEG_LOAD) begin
            if (soc_ctrl_i.new_eeg_data) begin
                /* cnt_7b_i holds current EEG data in patch
                   cnt_9b_i holds current patch */
                    IntResAddr_t addr = mem_map[EEG_INPUT_MEM] + IntResAddr_t'(int'(cnt_7b_i.cnt) + (int'(cnt_9b_i.cnt) << $clog2(PATCH_LEN)));
                    CompFx_t eeg_normalized = CompFx_t'({soc_ctrl_i.eeg, (Q_COMP-ADC_BITWIDTH)'(0)}); // Normalize to [0, 1]
                    write_int_res(addr, eeg_normalized, int_res_width[EEG_WIDTH], int_res_format[EEG_FORMAT]);
                    if (int'(cnt_7b_i.cnt) == PATCH_LEN-1) begin
                        cnt_7b_i.rst_n <= 1'b0;
                        if (int'(cnt_9b_i.cnt) == NUM_PATCHES-1) cnt_9b_i.rst_n <= 1'b0;
                        else cnt_9b_i.inc <= 1'b1;
                    end else cnt_7b_i.inc <= 1'b1;
            end
        end else if (cim_state == INFERENCE_RUNNING) begin
            unique case (current_inf_step)
                PATCH_PROJ_STEP: begin
                    /* cnt_7b_i holds current parameters row
                       cnt_9b_i holds current patch */

                    if ((mac_io.done || (cnt_7b_i.cnt == 0 && ~mac_io.busy)) && (int'(cnt_7b_i.cnt) != EMB_DEPTH-1)) begin
                        IntResAddr_t patch_addr = mem_map[EEG_INPUT_MEM] + IntResAddr_t'(int'(cnt_9b_i.cnt) << $clog2(EMB_DEPTH));
                        ParamAddr_t param_addr  = param_addr_map[PATCH_PROJ_KERNEL_PARAMS] + ParamAddr_t'(int'(cnt_7b_i.cnt) << $clog2(EMB_DEPTH));
                        ParamAddr_t bias_addr   = param_addr_map_bias[PATCH_PROJ_BIAS] + ParamAddr_t'(cnt_7b_i.cnt);
                        start_mac(patch_addr, IntResAddr_t'(param_addr), bias_addr, MODEL_PARAM, LINEAR_ACTIVATION, VectorLen_t'(PATCH_LEN), int_res_format[EEG_FORMAT],
                                  int_res_width[EEG_WIDTH], params_format[PATCH_PROJ_PARAM_FORMAT]);
                    end

                    if (mac_io.done) begin
                        IntResAddr_t int_res_write_addr = mem_map[PATCH_MEM] + IntResAddr_t'(int'(cnt_7b_i.cnt) + int'(cnt_9b_i.cnt) << $clog2(PATCH_LEN)); // Left shift instead of multiply since PATCH_LEN is a power of 2
                        write_int_res(int_res_write_addr, mac_io.out, int_res_width[PATCH_PROJ_OUTPUT_WIDTH], int_res_format[PATCH_PROJ_OUTPUT_FORMAT]);

                        // Update index control
                        if (int'(cnt_7b_i.cnt) == EMB_DEPTH-1) begin
                            cnt_7b_i.rst_n <= 1'b0;
                            if (int'(cnt_9b_i.cnt) == NUM_PATCHES-1) begin
                                cnt_9b_i.rst_n <= 1'b0;
                                current_inf_step <= CLASS_TOKEN_CONCAT_STEP;
                            end else cnt_9b_i.inc <= 1'b1;
                        end else cnt_7b_i.inc <= 1'b1;
                    end
                end
                CLASS_TOKEN_CONCAT_STEP: begin
                    cnt_7b_i.inc <= 1'b1;
                    delay_line_2b[0] <= cnt_7b_i.inc; // One cycle delay
                    cnt_9b_i.inc <= delay_line_2b[0];
                    if (int'(cnt_9b_i.cnt) == EMB_DEPTH) begin
                        delay_line_2b <= 'b0;
                        cnt_7b_i.rst_n <= 1'b0;
                        cnt_9b_i.rst_n <= 1'b0;
                        current_inf_step <= POS_EMB_STEP;
                    end else begin
                        ParamAddr_t read_addr = param_addr_map_bias[CLASS_TOKEN] + ParamAddr_t'(cnt_7b_i.cnt);
                        IntResAddr_t write_addr = mem_map[CLASS_TOKEN_MEM] + IntResAddr_t'(cnt_9b_i.cnt);
                        if (cnt_7b_i.inc) read_params(read_addr, params_format[CLASS_EMB_TOKEN_PARAM_FORMAT]);
                        if (cnt_9b_i.inc) write_int_res(write_addr, param_read_i.data, int_res_width[CLASS_EMB_TOKEN_WIDTH], int_res_format[CLASS_EMB_TOKEN_FORMAT]);
                    end
                end
                POS_EMB_STEP: begin
                    /* gen_cnt_7b holds the column
                    gen_cnt_9b holds the row */

                    // TODO: The variables are updated with blocking operators. They would be synthesized with non-blocking operators, so does int_res_addr_write need to be updated in a line before int_res_addr_read?

                    ParamAddr_t params_addr = param_addr_map[POS_EMB_PARAMS] + ParamAddr_t'(cnt_7b_i.cnt) + ParamAddr_t'(EMB_DEPTH*cnt_9b_i.cnt);
                    IntResAddr_t int_res_addr_read = mem_map[CLASS_TOKEN_MEM] + IntResAddr_t'(cnt_7b_i.cnt) + IntResAddr_t'(EMB_DEPTH*cnt_9b_i.cnt);
                    IntResAddr_t int_res_addr_write = int_res_addr_read - (mem_map[CLASS_TOKEN_MEM] - mem_map[POS_EMB_MEM]) - IntResAddr_t'('d4);

                    // Read
                    if (cnt_7b_i.inc) read_params(params_addr, params_format[POS_EMB_PARAM_FORMAT]);
                    if (cnt_7b_i.inc) read_int_res(int_res_addr_read, int_res_width[CLASS_EMB_TOKEN_WIDTH], int_res_format[CLASS_EMB_TOKEN_FORMAT]);

                    // Add
                    if (delay_line_2b[1]) start_add(param_read_i.data, int_res_read_i.data);

                    // Write
                    if (add_io_cim.done) write_int_res(int_res_addr_write, add_io_cim.out, int_res_width[POS_EMB_WIDTH], int_res_format[POS_EMB_FORMAT]);

                    // Counter control
                    cnt_7b_i.inc <= 1'b1;
                    delay_line_2b[0] <= param_read_cim_i.en;
                    delay_line_2b[1] <= delay_line_2b[0]; // One cycle delay
                    if (int'(cnt_7b_i.cnt) == EMB_DEPTH-2) begin
                        cnt_7b_i.rst_n <= 1'b0;
                        cnt_9b_i.inc <= 1'b1;
                    end

                    // Done
                    if (int_res_addr_write == IntResAddr_t'(int'(mem_map[POS_EMB_MEM]) + EMB_DEPTH*(NUM_PATCHES+1) - 1)) begin
                        current_inf_step <= ENC_LAYERNORM_1_1ST_HALF_STEP;
                        delay_line_2b <= 'b0;
                        cnt_7b_i.rst_n <= 1'b0;
                        cnt_9b_i.rst_n <= 1'b0;
                    end
                end
                ENC_LAYERNORM_1_1ST_HALF_STEP: begin
                    if ((ln_io.done || (cnt_7b_i.cnt == 0 && ~ln_io.busy)) && ~ln_io.start && (int'(cnt_7b_i.cnt) != NUM_PATCHES+1)) begin
                        IntResAddr_t input_starting_addr = mem_map[POS_EMB_MEM] + IntResAddr_t'(EMB_DEPTH*cnt_7b_i.cnt);
                        IntResAddr_t output_starting_addr = mem_map[ENC_LN1_MEM] + IntResAddr_t'(EMB_DEPTH*cnt_7b_i.cnt);
                        start_layernorm(FIRST_HALF, input_starting_addr, output_starting_addr, param_addr_map_bias[ENC_LAYERNORM_1_BETA], param_addr_map_bias[ENC_LAYERNORM_1_GAMMA],
                                        int_res_width[LN_INPUT_WIDTH], int_res_format[LN_INPUT_FORMAT], int_res_width[LN_OUTPUT_WIDTH],
                                        int_res_format[LN_OUTPUT_FORMAT], params_format[LN_PARAM_FORMAT]);
                    end

                    cnt_7b_i.inc <= ln_io.start;

                    if (ln_io.done && (int'(cnt_7b_i.cnt) == NUM_PATCHES+1)) begin
                        cnt_7b_i.rst_n <= 1'b0;
                        current_inf_step <= ENC_LAYERNORM_1_2ND_HALF_STEP;
                    end
                end
                default: begin
                end
            endcase
        end
    end

    // ----- MUX -----//
    always_comb begin : param_mem_MUX // TODO: Why does it claim that no latch is inferred if I use always_latch?
        // Write (only testbench writes to params)
        param_write_i.data_width = SINGLE_WIDTH;
        param_write_i.chip_en = 1'b1;
        param_write_i.en = param_write_tb_i.en;
        param_write_i.addr = param_write_tb_i.addr;
        param_write_i.data = param_write_tb_i.data;
        param_write_i.format = param_write_tb_i.format;

        // Read
        param_read_i.data_width = SINGLE_WIDTH;
        param_read_i.en = param_read_mac_i.en | param_read_cim_i.en | param_read_ln_i.en;
        param_read_mac_i.data = param_read_i.data;
        param_read_ln_i.data = param_read_i.data;
        if (param_read_mac_i.en) begin // MAC
            param_read_i.addr = param_read_mac_i.addr;
            param_read_i.format = param_read_mac_i.format;
        end else if (param_read_cim_i.en) begin
            param_read_i.addr = param_read_cim_i.addr;
            param_read_i.format = param_read_cim_i.format;
        end else if (param_read_ln_i.en) begin
            param_read_i.addr = param_read_ln_i.addr;
            param_read_i.format = param_read_ln_i.format;
        end
    end

    always_latch begin : int_res_mem_MUX
        // Write
        int_res_write_i.chip_en = 1'b1;
        int_res_write_i.en = int_res_write_tb_i.en | int_res_write_cim_i.en | int_res_write_ln_i.en;
        if (int_res_write_tb_i.en) begin
            int_res_write_i.addr = int_res_write_tb_i.addr;
            int_res_write_i.data = int_res_write_tb_i.data;
            int_res_write_i.format = int_res_write_tb_i.format;
            int_res_write_i.data_width = int_res_write_tb_i.data_width;
        end else if (int_res_write_cim_i.en) begin
            int_res_write_i.addr = int_res_write_cim_i.addr;
            int_res_write_i.data = int_res_write_cim_i.data;
            int_res_write_i.format = int_res_write_cim_i.format;
            int_res_write_i.data_width = int_res_write_cim_i.data_width;
        end else if (int_res_write_ln_i.en) begin
            int_res_write_i.addr = int_res_write_ln_i.addr;
            int_res_write_i.data = int_res_write_ln_i.data;
            int_res_write_i.format = int_res_write_ln_i.format;
            int_res_write_i.data_width = int_res_write_ln_i.data_width;
        end

        // Read
        int_res_read_i.en = int_res_read_mac_i.en | int_res_read_cim_i.en | int_res_read_ln_i.en;
        int_res_read_mac_i.data = int_res_read_i.data;
        int_res_read_cim_i.data = int_res_read_i.data;
        int_res_read_ln_i.data = int_res_read_i.data;
        if (int_res_read_mac_i.en) begin // MAC
            int_res_read_i.addr = int_res_read_mac_i.addr;
            int_res_read_i.data_width = int_res_read_mac_i.data_width;
            int_res_read_i.format = int_res_read_mac_i.format;
        end else if (int_res_read_cim_i.en) begin
            int_res_read_i.addr = int_res_read_cim_i.addr;
            int_res_read_i.data_width = int_res_read_cim_i.data_width;
            int_res_read_i.format = int_res_read_cim_i.format;
        end else if (int_res_read_ln_i.en) begin
            int_res_read_i.addr = int_res_read_ln_i.addr;
            int_res_read_i.data_width = int_res_read_ln_i.data_width;
            int_res_read_i.format = int_res_read_ln_i.format;
        end
    end

    always_latch begin : add_io_MUX
        if (add_io_exp.start) begin
            add_io.in_1 = add_io_exp.in_1;
            add_io.in_2 = add_io_exp.in_2;
        end else if (add_io_mac.start) begin
            add_io.in_1 = add_io_mac.in_1;
            add_io.in_2 = add_io_mac.in_2;
        end else if (add_io_cim.start) begin
            add_io.in_1 = add_io_cim.in_1;
            add_io.in_2 = add_io_cim.in_2;
        end else if (add_io_ln.start) begin
            add_io.in_1 = add_io_ln.in_1;
            add_io.in_2 = add_io_ln.in_2;
        end

        add_io.start = add_io_exp.start | add_io_mac.start | add_io_cim.start | add_io_ln.start;
        add_io_exp.out = add_io.out;
        add_io_exp.done = add_io.done;
        add_io_mac.out = add_io.out;
        add_io_mac.done = add_io.done;
        add_io_cim.out = add_io.out;
        add_io_cim.done = add_io.done;
        add_io_ln.out = add_io.out;
        add_io_ln.done = add_io.done;
    end

    always_latch begin : mult_io_MUX
        if (mult_io_exp.start) begin
            mult_io.in_1 = mult_io_exp.in_1;
            mult_io.in_2 = mult_io_exp.in_2;
        end else if (mult_io_mac.start) begin
            mult_io.in_1 = mult_io_mac.in_1;
            mult_io.in_2 = mult_io_mac.in_2;
        end else if (mult_io_ln.start) begin
            mult_io.in_1 = mult_io_ln.in_1;
            mult_io.in_2 = mult_io_ln.in_2;
        end

        mult_io.start = mult_io_exp.start | mult_io_mac.start | mult_io_ln.start;
        mult_io_exp.out = mult_io.out;
        mult_io_exp.done = mult_io.done;
        mult_io_mac.out = mult_io.out;
        mult_io_mac.done = mult_io.done;
        mult_io_ln.out = mult_io.out;
        mult_io_ln.done = mult_io.done;
    end

    always_latch begin : div_io_MUX
        if (div_io_mac.start) begin
            div_io.in_1 = div_io_mac.in_1;
            div_io.in_2 = div_io_mac.in_2;
        end else if (div_io_ln.start) begin
            div_io.in_1 = div_io_ln.in_1;
            div_io.in_2 = div_io_ln.in_2;
        end

        div_io.start = div_io_mac.start | div_io_ln.start;
        div_io_mac.out = div_io.out;
        div_io_mac.busy = div_io.busy;
        div_io_mac.done = div_io.done;
        div_io_ln.out = div_io.out;
        div_io_ln.busy = div_io.busy;
        div_io_ln.done = div_io.done;
    end

    always_latch begin : exp_io_MUX
        if (exp_io_mac.start) begin
            exp_io.in_1 = exp_io_mac.in_1;
        end

        exp_io.in_2 = CompFx_t'(0);
        exp_io.start = exp_io_mac.start;
        exp_io_mac.out = exp_io.out;
        exp_io_mac.busy = exp_io.busy;
        exp_io_mac.done = exp_io.done;
    end

    // ----- TASKS ----- //
    task automatic set_default_values();
        // Sets the default value for signals that do not persist cycle-to-cycle
        cnt_4b_i.inc <= 1'b0;
        cnt_7b_i.inc <= 1'b0;
        cnt_9b_i.inc <= 1'b0;
        cnt_4b_i.rst_n <= 1'b1;
        cnt_7b_i.rst_n <= 1'b1;
        cnt_9b_i.rst_n <= 1'b1;

        param_read_cim_i.en <= 1'b0;
        int_res_read_cim_i.en <= 1'b0;
        int_res_write_cim_i.en <= 1'b0;

        mac_io.start <= 1'b0;
        add_io_cim.start <= 1'b0;
        ln_io.start <= 1'b0;
    endtask

    task automatic reset();
        cim_state <= IDLE_CIM;
        current_inf_step <= PATCH_PROJ_STEP;

        cnt_4b_i.inc <= 1'b0;
        cnt_7b_i.inc <= 1'b0;
        cnt_9b_i.inc <= 1'b0;
        cnt_4b_i.rst_n <= 1'b0;
        cnt_7b_i.rst_n <= 1'b0;
        cnt_9b_i.rst_n <= 1'b0;

        mac_io.start <= 1'b0;
        add_io_cim.start <= 1'b0;
    endtask

    task write_int_res(input IntResAddr_t addr, input CompFx_t data, input DataWidth_t width, input FxFormatIntRes_t int_res_format);
        int_res_write_cim_i.en <= 1'b1;
        int_res_write_cim_i.addr <= addr;
        int_res_write_cim_i.data <= data;
        int_res_write_cim_i.data_width <= width;
        int_res_write_cim_i.format <= int_res_format;
    endtask

    task read_params(input ParamAddr_t addr, input FxFormatParams_t format);
        param_read_cim_i.en <= 1'b1;
        param_read_cim_i.addr <= addr;
        param_read_cim_i.format <= format;
    endtask

    task read_int_res(input IntResAddr_t addr, input DataWidth_t width, input FxFormatIntRes_t int_res_format);
        int_res_read_cim_i.en <= 1'b1;
        int_res_read_cim_i.addr <= addr;
        int_res_read_cim_i.data_width <= width;
        int_res_read_cim_i.format <= int_res_format;
    endtask

    task start_mac(input IntResAddr_t addr_1, input IntResAddr_t addr_2, input ParamAddr_t bias_addr, input ParamType_t param_type, input Activation_t act, input VectorLen_t len, input FxFormatIntRes_t int_res_input_format, input DataWidth_t int_res_read_width, input FxFormatParams_t params_read_format);
        mac_io.start <= 1'b1;
        mac_io_extra.start_addr_1 <= addr_1;
        mac_io_extra.start_addr_2 <= addr_2;
        mac_io_extra.param_type <= param_type;
        mac_io_extra.activation <= act;
        mac_io_extra.len <= len;
        mac_io_extra.bias_addr <= bias_addr;
        mac_casts_i.int_res_read_format <= int_res_input_format;
        mac_casts_i.int_res_read_width <= int_res_read_width;
        mac_casts_i.params_read_format <= params_read_format;
    endtask

    task start_add(CompFx_t in_1, CompFx_t in_2);
        add_io_cim.start <= 1'b1;
        add_io_cim.in_1 <= in_1;
        add_io_cim.in_2 <= in_2;
    endtask

    task start_layernorm(input HalfSelect_t half_select, input IntResAddr_t input_starting_addr, input IntResAddr_t output_starting_addr, input ParamAddr_t beta_addr, input ParamAddr_t gamma_addr, input DataWidth_t input_width, input FxFormatIntRes_t input_format, input DataWidth_t output_width, input FxFormatIntRes_t output_format, input FxFormatParams_t param_format);
        ln_io.start <= 1'b1;
        ln_io_extra.half_select <= half_select;
        ln_io_extra.start_addr_1 <= input_starting_addr;
        ln_io_extra.start_addr_2 <= output_starting_addr;
        ln_io_extra.start_addr_3 <= IntResAddr_t'(beta_addr);
        ln_io_extra.start_addr_4 <= IntResAddr_t'(gamma_addr);
        ln_casts_i.int_res_read_format <= input_format;
        ln_casts_i.int_res_write_format <= output_format;
        ln_casts_i.int_res_read_width <= input_width;
        ln_casts_i.int_res_write_width <= output_width;
        ln_casts_i.params_read_format <= param_format;
    endtask

    // ----- ASSERTIONS ----- //
    always_ff @ (posedge clk) begin : compute_mux_assertions
        assert (~(int_res_write_tb_i.en & int_res_write_cim_i.en & int_res_write_ln_i.en)) else $fatal("More than one source are trying to write to intermediate result memory simulatenously!");
        assert (~(int_res_read_cim_i.en & int_res_read_mac_i.en & int_res_read_ln_i.en)) else $fatal("More than one source are trying to read from intermediate results memory simulatenously!");
        assert (~(param_read_cim_i.en & param_read_mac_i.en & param_read_ln_i.en)) else $fatal("More than one source are trying to read from parameters result memory simulatenously!");

        assert (~(add_io_exp.start & add_io_mac.start & add_io_cim.start & add_io_ln.start)) else $fatal("More than one source are trying to start an add!");
        assert (~(mult_io_exp.start & mult_io_mac.start & mult_io_ln.start)) else $fatal("More than one source are trying to start a mult!");
        assert (~(div_io_mac.start & div_io_ln.start)) else $fatal("More than one source are trying to start a div!");
        assert (~(exp_io_mac.start & 0)) else $fatal("More than one source are trying to start an exp!");
    end
endmodule

`endif // _cim_centralized_vh_
