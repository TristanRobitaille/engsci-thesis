module cim_centralized #(
    parameter STANDALONE_TB = 0
)(
    input wire clk, rst
);

endmodule