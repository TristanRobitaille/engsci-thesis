`ifndef _master_vh_
`define _master_vh_

/*----- ENUM -----*/
    typedef enum logic [2:0] {
        MASTER_STATE_IDLE,
        MASTER_STATE_PARAM_LOAD,
        MASTER_STATE_SIGNAL_LOAD,
        MASTER_STATE_INFERENCE_RUNNING,
        MASTER_STATE_BROADCAST_MANAGEMENT,
        MASTER_STATE_WAITING_FOR_CIM_COMPLETION
    } MASTER_STATE_T;

    typedef enum logic [4:0] {
        PRE_LAYERNORM_1_TRANS_STEP,
        INTRA_LAYERNORM_1_TRANS_STEP,
        POST_LAYERNORM_1_TRANS_STEP,
        ENC_MHSA_DENSE_STEP,
        ENC_MHSA_Q_TRANS_STEP,
        ENC_MHSA_K_TRANS_STEP,
        ENC_MHSA_QK_T_STEP,
        ENC_MHSA_PRE_SOFTMAX_TRANS_STEP,
        ENC_MHSA_SOFTMAX_STEP,
        ENC_MHSA_V_MULT_STEP,
        ENC_MHSA_POST_V_TRANS_STEP,
        ENC_MHSA_POST_V_DENSE_STEP,
        PRE_LAYERNORM_2_TRANS_STEP,
        INTRA_LAYERNORM_2_TRANS_STEP,
        ENC_PRE_MLP_TRANSPOSE_STEP,
        ENC_MLP_DENSE_1_STEP,
        ENC_MLP_DENSE_2_TRANSPOSE_STEP,
        ENC_MLP_DENSE_2_AND_SUM_STEP,
        PRE_LAYERNORM_3_TRANS_STEP,
        INTRA_LAYERNORM_3_TRANS_STEP,
        PRE_MLP_HEAD_DENSE_TRANS_STEP,
        MLP_HEAD_DENSE_1_STEP,
        PRE_MLP_HEAD_DENSE_2_TRANS_STEP,
        MLP_HEAD_DENSE_2_STEP,
        MLP_HEAD_SOFTMAX_TRANS_STEP,
        SOFTMAX_AVERAGING,
        INFERENCE_FINISHED
    } HIGH_LEVEL_INFERENCE_STEP_T;

`endif
