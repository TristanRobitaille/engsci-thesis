`ifndef _master_fcn_vh_
`define _master_fcn_vh_

`include "../types.svh"

/*----- FUNCTIONS -----*/
function automatic void param_to_send();
endfunction

`endif
